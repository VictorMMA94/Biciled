Library ieee;
Use ieee.std_logic_1164.all;
Use ieee.std_logic_unsigned.all;
Use IEEE.std_logic_arith.all;
Use work.mis_componentes.all;
---------------------------------------------------------------------------------------------------------
ENTITY SENALETICA_BICI IS
PORT(	START: 					In std_logic;
		LEFT_BUTTON: 			In std_logic;
		RIGHT_BUTTON: 			In std_logic;
		MOSTRAR_BUTTON: 		In std_logic;
		RESET: 					In std_logic;
		MANUAL_AUTO:			In std_logic;
		CLOCK_MANUAL: 			In std_logic;
		CLOCK_FPGA: 			In std_logic;
		CLOCK_1KHz:				In std_logic;
		LUCES_LEDS:				Out std_logic_vector(19 downto 0);
		DISPLAY_MIL:			Out std_logic_vector(6 downto 0);
		DISPLAY_CENTENAS:		Out std_logic_vector(6 downto 0);
		DISPLAY_DECENAS:		Out std_logic_vector(6 downto 0);
		DISPLAY_UNIDADES:		Out std_logic_vector(6 downto 0));
		
END SENALETICA_BICI; 
---------------------------------------------------------------------------------------------------------
ARCHITECTURE estructural OF SENALETICA_BICI IS
-------------------------------------------------------------------------------------------------------------

SIGNAL RL, RR, NORMAL, EMERGENCIA: std_logic;
SIGNAL LOAD_REG, RESET_REG, CAMBIA_USADO: std_logic;
SIGNAL LUCES_1, LUCES_2, LUCES_3, LUCES_4: std_logic_vector(19 downto 0);
SIGNAL S1, S0: std_logic;
SIGNAL RESET_1, CLOCK_1K: std_logic;
SIGNAL MILISEGUNDOS: std_logic_vector(8 downto 0);
SIGNAL CAMBIA: std_logic;
SIGNAL EN_TIME, RESET_TIME: std_logic;
SIGNAL CLOCK_USADO, CLOCK_USADO_CENT, CLOCK_DEC, CLOCK_CENT, CLOCK_MIL : std_logic;
SIGNAL UNIDADES, DECENAS, CENTENAS, MIL: std_logic_vector(3 downto 0);
SIGNAL FIN_SECUENCIA, PRENDE, EN_DISPLAY, RESET_FF: std_logic;
SIGNAL SIN_USO: std_logic;

-------------------------------------------------------------------------------------------------------------
BEGIN
	PROCESS(MILISEGUNDOS, MIL)
	BEGIN
	IF MILISEGUNDOS="111110100" THEN CAMBIA<='1'; ELSE CAMBIA<='0'; END IF;
	IF (MIL="0101" OR MIL>"0101") THEN FIN_SECUENCIA<='1'; ELSE FIN_SECUENCIA<='0'; END IF;
	END PROCESS;
	
	REGISTRO_DESPLAZAMIENTO_IZQUIERDA: registro_d_i PORT MAP(RESET_REG, CAMBIA_USADO OR LOAD_REG, RL OR LOAD_REG, LOAD_REG, "00000000000000000001", LUCES_1);
	REGISTRO_DESPLAZAMIENTO_DERECHA: registro_i_d PORT MAP(RESET_REG, CAMBIA_USADO OR LOAD_REG, RR OR LOAD_REG, LOAD_REG, "10000000000000000000", LUCES_2);
	REGISTRO_SOSTENIMIENYO_ALTERNADO: registro_alternado PORT MAP( RESET_REG, CAMBIA_USADO OR LOAD_REG, NORMAL, LOAD_REG, "11110000111100001111", LUCES_3);
	REGISTRO_SOSTENIMIENYO_ON_OFF: registro_ON_OFF PORT MAP( RESET_REG, CAMBIA_USADO OR LOAD_REG, EMERGENCIA OR LOAD_REG, LOAD_REG, "00000000000000000000", LUCES_4);
	MULTIPLEXADOR_4_A_1_LUCES: MUX_4to1 PORT MAP( LUCES_3, LUCES_2, LUCES_1, LUCES_4, LUCES_LEDS, S1&S0); 
	DEMULTIPLEXADOR_1_A_4_ENABLES_LUCES: DEMUX_4to1 PORT MAP( '1', NORMAL, RR, RL, EMERGENCIA, S1&S0);
	MULTIPLEXADOR_2_A_1_CAMBIADOR: MUX_2_1 PORT MAP( CAMBIA, CLOCK_MANUAL, MANUAL_AUTO, CAMBIA_USADO); 
	MULTIPLEXADOR_2_A_1_CLOCK_UNIDADES: MUX_2_1 PORT MAP( CLOCK_1KHz, '0', MANUAL_AUTO, CLOCK_USADO_CENT); 
	MULTIPLEXADOR_2_A_1_CLOCK_CENTENAS: MUX_2_1 PORT MAP( CLOCK_CENT, CLOCK_MANUAL, MANUAL_AUTO, CLOCK_USADO); 
	FLIP_FLOP_DISPLAY: FF_tipoD PORT MAP( '1', PRENDE, (RESET_FF OR FIN_SECUENCIA), PRENDE, EN_DISPLAY);
	CONTADOR_MILISEGUNDOS: CONTADOR_UP_0_500 PORT MAP(	RESET_1, CLOCK_1KHz, '1', '0', "000000000", MILISEGUNDOS);
	CONTADOR_TIME_UNIDADES: CONTADOR_UP_0TO9 PORT MAP(	EN_TIME, '0', RESET_TIME, CLOCK_USADO, "0000", CLOCK_DEC, UNIDADES);
	CONTADOR_TIME_DECENAS: CONTADOR_UP_0TO9 PORT MAP( EN_TIME, '0', RESET_TIME, CLOCK_DEC, "0000", CLOCK_CENT, DECENAS);
	CONTADOR_TIME_CENTENAS: CONTADOR_UP_0TO9 PORT MAP( EN_TIME, '0', RESET_TIME, CLOCK_USADO_CENT, "0000", CLOCK_MIL, CENTENAS);
	CONTADOR_TIME_MILES: CONTADOR_UP_0TO9 PORT MAP( EN_TIME, '0', RESET_TIME, CLOCK_MIL, "0000", SIN_USO, MIL);
	DISPLAY_7SEG_U: DECODER_7SEG PORT MAP ( UNIDADES, EN_DISPLAY, DISPLAY_UNIDADES);
	DISPLAY_7SEG_D: DECODER_7SEG PORT MAP ( DECENAS, EN_DISPLAY, DISPLAY_DECENAS);
	DISPLAY_7SEG_C: DECODER_7SEG PORT MAP ( CENTENAS, EN_DISPLAY, DISPLAY_CENTENAS);
	DISPLAY_7SEG_M: DECODER_7SEG PORT MAP ( MIL, EN_DISPLAY, DISPLAY_MIL);
	CONTROLADOR: CONTROLADORA_MSS PORT MAP( START, LEFT_BUTTON, RIGHT_BUTTON, MOSTRAR_BUTTON, FIN_SECUENCIA, RESET, CLOCK_FPGA, LOAD_REG, RESET_REG, S1, S0, RESET_1, EN_TIME, RESET_TIME, RESET_FF, PRENDE);
	
END estructural;